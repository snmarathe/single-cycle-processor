`include "instruction_memory.v"
`include "program_counter.v"
`include "increment_pc.v"
`include "registers.v"
`include "data_memory.v"
`include "ALU.v"
`include "ALU_ctrl.v"
`include "ALU_operand_mux.v"
`include "send_to_reg_mux.v"
`include "sign_extend.v"
`include "branch_addr.v"
`include "branch_mux.v"
`include "jump_addr.v"
`include "jump_mux.v"
`include "flags.v"

module processor(

);

endmodule
